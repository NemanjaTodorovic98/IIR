`ifndef IIR_SEQ_PKG_SV
 `define IIR_SEQ_PKG_SV
package iir_seq_pkg;
   import uvm_pkg::*;      // import the UVM library
 `include "uvm_macros.svh" // Include the UVM macros
  import iir_agent_pkg::iir_seq_item;
   import iir_agent_pkg::iir_sequencer;
 `include "iir_base_seq.sv"
 `include "iir_simple_seq.sv"
     endpackage 
`endif
