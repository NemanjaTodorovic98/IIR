library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package types is

     type logic_vector_array_type_fixed is array (0 to 19) of std_logic_vector(31 downto 0);

end package types;